package build_id is
constant BUILD_DATE : string := "230515";
constant BUILD_TIME : string := "181623";
end build_id;
